* ring_oscillator_3

.subckt ring_oscillator_3 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=1.0817986949047222 d_WP=1.0192112229511558 d_LN=1.0048554239402694 d_WN=1.0886572404937314 d_TOXEP=1.0555764851965357 d_TOXEN=1.055541521310898
x2 n1 n2 inverter d_LP=1.0001014777490156 d_WP=1.0620723184267356 d_LN=1.0190926333481856 d_WN=0.971640640305692 d_TOXEP=0.9826740202482269 d_TOXEN=1.0163748591924295
x3 n2 n3 inverter d_LP=1.0414134508621802 d_WP=0.9746312513279255 d_LN=1.069949334187812 d_WN=0.874031681137682 d_TOXEP=0.9655986981384593 d_TOXEN=1.0333814211571513
x4 n3 n4 inverter d_LP=0.9213597846613747 d_WP=0.9872686400749198 d_LN=1.031783472740848 d_WN=1.0464146618587193 d_TOXEP=0.961131349585467 d_TOXEN=1.0010388261820984
x5 n4 n5 inverter d_LP=0.9580988833181117 d_WP=1.033851694843311 d_LN=0.9130506841065653 d_WN=1.023996804419223 d_TOXEP=0.9756767970770881 d_TOXEN=1.0102339556228013
x6 n5 n6 inverter d_LP=0.8715383766400621 d_WP=0.9140287137501429 d_LN=1.0607277395197139 d_WN=1.0906081960159393 d_TOXEP=1.0103841280260564 d_TOXEN=0.977113407213474
x7 n6 n7 inverter d_LP=1.023558208100207 d_WP=1.0435373066196838 d_LN=0.8966898450139752 d_WN=1.0198609282600262 d_TOXEP=1.039018934860496 d_TOXEN=0.9661815541033497
x8 n7 n8 inverter d_LP=1.0738596143529318 d_WP=0.9181313911299456 d_LN=1.0847930884881862 d_WN=0.9274416486841941 d_TOXEP=0.9442566351748297 d_TOXEN=1.0650056256645655
x9 n8 n9 inverter d_LP=1.0860293154057128 d_WP=0.9625518780202634 d_LN=0.9815033053984183 d_WN=1.0408454322215064 d_TOXEP=1.0117841685948157 d_TOXEN=0.9252781850792499
x10 n9 n10 inverter d_LP=0.9287879563789726 d_WP=1.0572995158210177 d_LN=1.0761365750316507 d_WN=1.0830045461977804 d_TOXEP=0.9558974003233539 d_TOXEN=0.9822703772996177
x11 n10 n11 inverter d_LP=0.9912521344721491 d_WP=0.9569275272679276 d_LN=1.0566230981331544 d_WN=0.9823779596662636 d_TOXEP=0.9639802749933433 d_TOXEN=1.0124649894200655
x12 n11 n12 inverter d_LP=0.970501978231526 d_WP=0.9881477433255955 d_LN=0.9989806450099404 d_WN=0.9620009560264922 d_TOXEP=1.0727634839631002 d_TOXEN=0.9529398213781061
.ends ring_oscillator_3

