* ring_oscillator_1

.subckt ring_oscillator_1 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=1.01779547322775 d_WP=0.9670029164311269 d_LN=1.0157101180921944 d_WN=0.9978064261029738 d_TOXEP=1.0674893083937693 d_TOXEN=0.9772425232744327
x2 n1 n2 inverter d_LP=1.0830153280335655 d_WP=0.9434072211164056 d_LN=0.9418085090526195 d_WN=0.9664890116760175 d_TOXEP=0.9256948536110349 d_TOXEN=0.983805574154075
x3 n2 n3 inverter d_LP=1.0700289183820564 d_WP=1.1099134235272208 d_LN=0.8589943775060953 d_WN=0.8953688343472761 d_TOXEP=0.9187681991693262 d_TOXEN=0.9882159547126222
x4 n3 n4 inverter d_LP=1.0146399494557918 d_WP=0.9795147285680309 d_LN=0.9881311933892011 d_WN=1.0413273675388284 d_TOXEP=0.9481176960562487 d_TOXEN=1.0571059654274308
x5 n4 n5 inverter d_LP=1.031275585094544 d_WP=1.0133317209428048 d_LN=0.8988446233616939 d_WN=1.044417973572892 d_TOXEP=1.0498315650897603 d_TOXEN=0.9806783506547648
x6 n5 n6 inverter d_LP=1.0560997771107326 d_WP=1.0317650283702722 d_LN=0.9100078915312573 d_WN=1.0110172005973619 d_TOXEP=0.9263914702342599 d_TOXEN=1.0389531593028813
x7 n6 n7 inverter d_LP=0.9379393991739763 d_WP=0.9839605709951869 d_LN=0.9322082318326208 d_WN=1.0100236773686897 d_TOXEP=0.9589862222975726 d_TOXEN=0.9632932385652433
x8 n7 n8 inverter d_LP=1.1097236409399245 d_WP=1.0824679663953447 d_LN=0.9621068339341514 d_WN=0.9851082078398243 d_TOXEP=0.927256408121193 d_TOXEN=0.9180890374324376
x9 n8 n9 inverter d_LP=1.0051480346918455 d_WP=0.9481481613512754 d_LN=0.964767927116777 d_WN=1.0192124426983948 d_TOXEP=1.071696349689095 d_TOXEN=1.0523549951176436
x10 n9 n10 inverter d_LP=1.145712550777329 d_WP=1.1062625946629288 d_LN=1.1332111904203577 d_WN=1.0540023460257504 d_TOXEP=1.0246117247705855 d_TOXEN=0.9892555145550105
x11 n10 n11 inverter d_LP=0.9336737039036749 d_WP=1.1007506351346812 d_LN=1.0166016851649888 d_WN=1.0615060616833603 d_TOXEP=1.0082293422464979 d_TOXEN=1.0846447124246414
x12 n11 n12 inverter d_LP=1.0599372928227158 d_WP=0.9840433338828507 d_LN=1.0113560929534788 d_WN=1.0068574407860174 d_TOXEP=1.0078242499612653 d_TOXEN=1.0018977953189423
.ends ring_oscillator_1

