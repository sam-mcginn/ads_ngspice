* ring_oscillator_6

.subckt ring_oscillator_6 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=0.9880009573110958 d_WP=1.0654225916267093 d_LN=0.990565544562941 d_WN=1.047490447756488 d_TOXEP=0.9942379646159482 d_TOXEN=1.023821317529591
x2 n1 n2 inverter d_LP=0.9998757504001647 d_WP=1.0136498647841916 d_LN=0.9733321915812193 d_WN=0.8693465267038634 d_TOXEP=1.0075200770392592 d_TOXEN=1.0513511220112342
x3 n2 n3 inverter d_LP=1.0161094444341245 d_WP=1.1172282397300368 d_LN=0.9590555146933394 d_WN=1.010522548243045 d_TOXEP=1.0183202150724053 d_TOXEN=0.959317451446451
x4 n3 n4 inverter d_LP=1.0341605558569318 d_WP=1.0957338097944567 d_LN=1.0120430517518335 d_WN=1.0796146135465665 d_TOXEP=1.0459100364695002 d_TOXEN=0.9521226130356406
x5 n4 n5 inverter d_LP=1.072730605770769 d_WP=0.8899651482259068 d_LN=1.0657590480511259 d_WN=0.9959345921429313 d_TOXEP=0.9664287646699962 d_TOXEN=0.9926704982696404
x6 n5 n6 inverter d_LP=1.0197563244089438 d_WP=0.9702604175307176 d_LN=0.9070570905947073 d_WN=0.9160589200372852 d_TOXEP=1.0002721901852631 d_TOXEN=1.0219692641379439
x7 n6 n7 inverter d_LP=1.0356932934388898 d_WP=1.0724152941717988 d_LN=0.9232577917899036 d_WN=0.9987858560950641 d_TOXEP=1.0608136262934742 d_TOXEN=1.0107718133806687
x8 n7 n8 inverter d_LP=0.9947609550337557 d_WP=0.9928768640708088 d_LN=1.010395057525492 d_WN=0.9359326254697753 d_TOXEP=1.006616290320113 d_TOXEN=0.9878796281576157
x9 n8 n9 inverter d_LP=0.9968249026165558 d_WP=0.9745462290742569 d_LN=0.909416823653956 d_WN=1.0646780993691374 d_TOXEP=0.9667218515717715 d_TOXEN=1.0486679168299753
x10 n9 n10 inverter d_LP=1.0061749969051477 d_WP=1.076622687041177 d_LN=1.0522210705066553 d_WN=0.9270588877407552 d_TOXEP=1.0013085135442428 d_TOXEN=1.019021238640789
x11 n10 n11 inverter d_LP=1.0062544879889728 d_WP=0.9821850176329995 d_LN=1.0553082559911047 d_WN=0.9727739804746847 d_TOXEP=0.9415253897986229 d_TOXEN=0.9590355632833105
x12 n11 n12 inverter d_LP=1.0979709022461221 d_WP=0.9528982007085123 d_LN=1.0258307082018472 d_WN=1.018891196681955 d_TOXEP=1.0004418609758532 d_TOXEN=1.0388599722615481
.ends ring_oscillator_6

