* ring_oscillator_0
.subckt ring_oscillator_0 enable n12
.include nand2.sp
.include inverter.sp

x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=1.100573571207846 d_WP=1.082713055226178 d_LN=1.0648283345905833 d_WN=1.0037793410393163 d_TOXEP=0.9534063770484567 d_TOXEN=1.0201006777262773
x2 n1 n2 inverter d_LP=0.998174326434556 d_WP=1.0566650779995008 d_LN=0.9617222353476761 d_WN=1.0620597701892356 d_TOXEP=0.9433343487279644 d_TOXEN=1.0453184058550777
x3 n2 n3 inverter d_LP=0.9264719408535405 d_WP=1.0826548550889727 d_LN=1.099618972226955 d_WN=0.9112280321002052 d_TOXEP=1.0031528380101473 d_TOXEN=0.9873889442186708
x4 n3 n4 inverter d_LP=1.083868415376665 d_WP=0.9926350670859826 d_LN=0.9990043668975369 d_WN=1.0396642004205838 d_TOXEP=0.9797423977245088 d_TOXEN=0.9820286755098075
x5 n4 n5 inverter d_LP=1.0292149393708319 d_WP=0.9693877008442382 d_LN=1.1098203070993078 d_WN=0.9635635064113686 d_TOXEP=0.9671455003534595 d_TOXEN=0.9393797049913162
x6 n5 n6 inverter d_LP=0.9296362771326849 d_WP=0.997010706409818 d_LN=1.0846239768213566 d_WN=0.9362906622534354 d_TOXEP=1.0089388831031634 d_TOXEN=1.0556747978807504
x7 n6 n7 inverter d_LP=1.0359361009562542 d_WP=0.9142842329206413 d_LN=0.8668489733358969 d_WN=0.9043719056246878 d_TOXEP=0.9279394171457882 d_TOXEN=1.0170675524220991
x8 n7 n8 inverter d_LP=0.9070925423184608 d_WP=1.1163691506696838 d_LN=1.1150394605348664 d_WN=0.9566600776359057 d_TOXEP=0.9176055616240458 d_TOXEN=1.022619235008784
x9 n8 n9 inverter d_LP=1.0530815331780607 d_WP=1.063432147284455 d_LN=1.0533198096887595 d_WN=0.9744397696313025 d_TOXEP=0.9414884128584228 d_TOXEN=1.0307141784503444
x10 n9 n10 inverter d_LP=0.9770309299522976 d_WP=0.8773959259191124 d_LN=0.912080757593361 d_WN=0.9994539129449623 d_TOXEP=0.9798407346147173 d_TOXEN=0.9736739250305385
x11 n10 n11 inverter d_LP=1.0980420783644333 d_WP=1.1059556426449768 d_LN=0.9857617216518205 d_WN=0.9897936720537368 d_TOXEP=1.0455796390923846 d_TOXEN=1.0316475952387787
x12 n11 n12 inverter d_LP=0.9668758096976683 d_WP=1.061159316084019 d_LN=0.8825503410471582 d_WN=1.0051659496107404 d_TOXEP=0.9884265823166201 d_TOXEN=0.968628574249091
.ends ring_oscillator_0

