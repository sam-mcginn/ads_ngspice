* ring_oscillator_5

.subckt ring_oscillator_5 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=1.0204352844360847 d_WP=1.1159520133697474 d_LN=0.9386498841251916 d_WN=1.0992461305790397 d_TOXEP=0.998035656542776 d_TOXEN=0.9829191728773082
x2 n1 n2 inverter d_LP=0.889274325244059 d_WP=0.933982839765641 d_LN=0.9993049386820656 d_WN=0.9922433587568862 d_TOXEP=0.9182241707100831 d_TOXEN=1.0150970487242437
x3 n2 n3 inverter d_LP=1.0490534359601922 d_WP=0.9456159884448895 d_LN=0.9263417709289423 d_WN=1.0118607993213162 d_TOXEP=0.9227149191574153 d_TOXEN=1.0696284402294145
x4 n3 n4 inverter d_LP=0.9339965204173741 d_WP=0.9580279908776307 d_LN=1.0681689729078752 d_WN=1.0240866968423201 d_TOXEP=1.0219392592135546 d_TOXEN=0.9839424936628295
x5 n4 n5 inverter d_LP=1.1064000500355398 d_WP=0.9596109271345349 d_LN=1.0527963238401299 d_WN=0.8829696852369018 d_TOXEP=0.9517103155190122 d_TOXEN=1.0095084798284066
x6 n5 n6 inverter d_LP=1.0318461058320638 d_WP=0.9405311850620386 d_LN=0.9821432588105729 d_WN=0.9512301781898335 d_TOXEP=0.9666020879764455 d_TOXEN=1.0326824446207805
x7 n6 n7 inverter d_LP=1.0242432102786734 d_WP=0.9324492596725568 d_LN=0.9970955188135162 d_WN=1.0257844068306874 d_TOXEP=0.9427217523506823 d_TOXEN=1.028386450897552
x8 n7 n8 inverter d_LP=1.0576950661609477 d_WP=1.0495409944551506 d_LN=0.9088196453082211 d_WN=1.0568740446567866 d_TOXEP=0.9648031943826976 d_TOXEN=1.0280849382365214
x9 n8 n9 inverter d_LP=1.1378182592292747 d_WP=1.0249258306025928 d_LN=0.9913802781083491 d_WN=0.91552344704904 d_TOXEP=1.0139968942447868 d_TOXEN=0.9823708552138656
x10 n9 n10 inverter d_LP=0.9873368164890547 d_WP=0.8968869915326577 d_LN=1.0254516050666511 d_WN=0.8756245588421906 d_TOXEP=1.020189136552214 d_TOXEN=0.99574074119529
x11 n10 n11 inverter d_LP=0.8716000180687528 d_WP=1.0044800947685928 d_LN=0.8666946527116683 d_WN=1.0468918579329927 d_TOXEP=0.9533606434283461 d_TOXEN=0.9859821699880343
x12 n11 n12 inverter d_LP=0.9258430124699724 d_WP=0.9062885457095307 d_LN=0.9726460049009723 d_WN=1.0190468406268813 d_TOXEP=1.0313226957892403 d_TOXEN=0.9840288457085961
.ends ring_oscillator_5

