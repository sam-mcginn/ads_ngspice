* ring_oscillator_7

.subckt ring_oscillator_7 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=0.9771520945823814 d_WP=0.9574488681700692 d_LN=0.9357986207561174 d_WN=1.0081154686174165 d_TOXEP=0.9013463607664131 d_TOXEN=0.9266914692333523
x2 n1 n2 inverter d_LP=1.0079797802644699 d_WP=0.9874285677536425 d_LN=0.9783389725851391 d_WN=0.9978010172271998 d_TOXEP=0.9544654223894355 d_TOXEN=0.9858918468356006
x3 n2 n3 inverter d_LP=1.0016642192092666 d_WP=0.9874523811201656 d_LN=0.9693893113805435 d_WN=1.0372770516154726 d_TOXEP=0.9924044602726846 d_TOXEN=1.0338510680268376
x4 n3 n4 inverter d_LP=1.118416229445725 d_WP=1.0083637312949574 d_LN=1.016176931238204 d_WN=0.9845804307022368 d_TOXEP=1.010743429165481 d_TOXEN=0.9901206481810364
x5 n4 n5 inverter d_LP=0.9473444176441959 d_WP=1.029902900553985 d_LN=1.062090480974866 d_WN=0.9628825604126099 d_TOXEP=1.0155067623798 d_TOXEN=0.9979225723683971
x6 n5 n6 inverter d_LP=1.0759779966625391 d_WP=1.071074480916122 d_LN=1.0043317164172236 d_WN=1.0062592248422504 d_TOXEP=1.0369159761126607 d_TOXEN=1.061539551045091
x7 n6 n7 inverter d_LP=1.0343889347664004 d_WP=1.0502279302334157 d_LN=1.109152110045906 d_WN=1.0202241354391504 d_TOXEP=0.9871744165874188 d_TOXEN=1.0318648644308541
x8 n7 n8 inverter d_LP=1.1155007114384066 d_WP=0.9599774157383176 d_LN=0.9355731658006012 d_WN=1.0263599287230736 d_TOXEP=1.0652225496282484 d_TOXEN=0.9972920225509041
x9 n8 n9 inverter d_LP=0.925058496312847 d_WP=0.9249425401236955 d_LN=0.9175772477939241 d_WN=0.9803984468857405 d_TOXEP=1.0165144945630273 d_TOXEN=0.9744580494778826
x10 n9 n10 inverter d_LP=0.9623802897913566 d_WP=1.0624284556810564 d_LN=0.9976079233613239 d_WN=0.9388070785881316 d_TOXEP=1.0351122004940734 d_TOXEN=1.0730950505257677
x11 n10 n11 inverter d_LP=0.9205295425513936 d_WP=0.9517879161751527 d_LN=1.0263020511257535 d_WN=0.9594215657291427 d_TOXEP=1.030552617449172 d_TOXEN=0.9360645171364999
x12 n11 n12 inverter d_LP=0.9137803491936031 d_WP=0.9381280694143156 d_LN=1.0252021646307607 d_WN=0.9896656751383004 d_TOXEP=1.0222432889316326 d_TOXEN=1.002239953793119
.ends ring_oscillator_7

