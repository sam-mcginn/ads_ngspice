* ring_oscillator_2

.subckt ring_oscillator_2 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=0.9555893723279358 d_WP=0.933564810270283 d_LN=1.0639480291865568 d_WN=0.9741853748991264 d_TOXEP=0.9511274529650514 d_TOXEN=0.9579698336905095
x2 n1 n2 inverter d_LP=0.9761894678808364 d_WP=0.980996665518905 d_LN=0.9659681729414948 d_WN=0.9793756372292344 d_TOXEP=1.0169254484666885 d_TOXEN=0.9788344404552947
x3 n2 n3 inverter d_LP=0.9543196591693639 d_WP=0.9294647699257981 d_LN=0.8529608531505927 d_WN=1.049206184719142 d_TOXEP=0.9314118233018447 d_TOXEN=0.9627338647491259
x4 n3 n4 inverter d_LP=0.9704670038524754 d_WP=1.0004138636643862 d_LN=1.0456470321143079 d_WN=0.9854961559301532 d_TOXEP=0.9299608623767546 d_TOXEN=1.0254363281170118
x5 n4 n5 inverter d_LP=1.1489369016713162 d_WP=0.9972116197423734 d_LN=1.0937079197943476 d_WN=0.9710702144946949 d_TOXEP=1.0818370547509986 d_TOXEN=1.0094067889603011
x6 n5 n6 inverter d_LP=1.0987214378248056 d_WP=1.1432227515767968 d_LN=1.02308161610236 d_WN=0.9950011095377351 d_TOXEP=1.049556721720676 d_TOXEN=0.9181356191845395
x7 n6 n7 inverter d_LP=1.0386777846531001 d_WP=1.0629494536894863 d_LN=1.0206348083802244 d_WN=0.9594485013969231 d_TOXEP=1.0234229405543218 d_TOXEN=0.958305252050862
x8 n7 n8 inverter d_LP=0.9790635134184382 d_WP=1.0216302226475307 d_LN=0.928045901699226 d_WN=0.9925120272127865 d_TOXEP=1.0262120920009055 d_TOXEN=1.0565511230349482
x9 n8 n9 inverter d_LP=1.0700182743644264 d_WP=0.9462278496680481 d_LN=1.0652410251910045 d_WN=0.9545474189528917 d_TOXEP=0.9383107906475885 d_TOXEN=1.0296607939833695
x10 n9 n10 inverter d_LP=0.9182064334098982 d_WP=0.9593830504659187 d_LN=1.0202442235477178 d_WN=1.1377830098110238 d_TOXEP=0.9323038100391285 d_TOXEN=0.9481341533919405
x11 n10 n11 inverter d_LP=1.008711968179581 d_WP=1.0545259052013856 d_LN=1.0213031160422952 d_WN=1.079244955393782 d_TOXEP=0.9378684065517059 d_TOXEN=0.9590002250278093
x12 n11 n12 inverter d_LP=1.0332509998611565 d_WP=0.9153960028621974 d_LN=0.9485044353375751 d_WN=0.9799350556612112 d_TOXEP=0.9029657064276133 d_TOXEN=0.9957456944795082
.ends ring_oscillator_2

