* ring_oscillator_4
.subckt ring_oscillator_4 enable n12
.include nand2.sp
.include inverter.sp
x0 enable n12 n0 nand2
x1 n0 n1 inverter d_LP=1.0034183137997632 d_WP=1.0120710417902525 d_LN=1.0666316525357906 d_WN=0.859567141766236 d_TOXEP=1.0250902467704093 d_TOXEN=1.014401980305568
x2 n1 n2 inverter d_LP=1.081741331421806 d_WP=1.1196830145742533 d_LN=1.1032750333215608 d_WN=1.0845273471603696 d_TOXEP=0.910469259421341 d_TOXEN=1.0030192231079318
x3 n2 n3 inverter d_LP=1.0049036844753907 d_WP=0.976504365102244 d_LN=1.0310354208211279 d_WN=1.0174722717943887 d_TOXEP=1.0600418531969873 d_TOXEN=0.9909434026754903
x4 n3 n4 inverter d_LP=1.0097600524400823 d_WP=0.9462571278358901 d_LN=1.0558846869570717 d_WN=1.128259273540142 d_TOXEP=1.0062944155377271 d_TOXEN=1.0793867522786733
x5 n4 n5 inverter d_LP=1.035043354113221 d_WP=1.0563558440992482 d_LN=0.8930498838850012 d_WN=0.9249186869280405 d_TOXEP=1.003629427663011 d_TOXEN=1.0445667286285503
x6 n5 n6 inverter d_LP=0.9709984076911776 d_WP=1.0362393160812338 d_LN=0.9997520586672668 d_WN=1.007487190456185 d_TOXEP=0.9500423549900324 d_TOXEN=1.0884003302960104
x7 n6 n7 inverter d_LP=0.9270070614875308 d_WP=0.9276083802901454 d_LN=0.9154543108717883 d_WN=0.9088580546473484 d_TOXEP=0.9851011097594751 d_TOXEN=1.0228960567970107
x8 n7 n8 inverter d_LP=1.104730397087546 d_WP=1.0219806364419328 d_LN=1.1024186124882323 d_WN=0.9368194075904259 d_TOXEP=1.0217293123296236 d_TOXEN=1.0007385749629376
x9 n8 n9 inverter d_LP=0.9032198399247329 d_WP=1.0211371598934316 d_LN=1.03645384139508 d_WN=0.9485236733105855 d_TOXEP=1.0903033299611287 d_TOXEN=0.999905829797339
x10 n9 n10 inverter d_LP=0.9041833897444845 d_WP=1.0234039424906365 d_LN=0.9366583502822576 d_WN=1.0078733070779773 d_TOXEP=1.0173517620976533 d_TOXEN=0.9851467119110271
x11 n10 n11 inverter d_LP=1.005343389476217 d_WP=0.9393756804155718 d_LN=1.0200650275937884 d_WN=1.0930905507416693 d_TOXEP=0.9648730020416608 d_TOXEN=1.0237409166770615
x12 n11 n12 inverter d_LP=1.0531369885827198 d_WP=0.9945770540473909 d_LN=0.9488744205055349 d_WN=0.9775066599205671 d_TOXEP=1.0160603358899967 d_TOXEN=0.9930708581752515
.ends ring_oscillator_4

